
// DEFINES 
`define __FILE__ "NA.v"
`define __LINE__ 0
`define DVT_PATCH

// CONFIGURATION FILES (libmap) 
`include "/home/student/akamien/VDIC/Lab0/apple.sv"
`include "/home/student/akamien/VDIC/Lab0/apple_tb.sv"
