
// DEFINES 
`define __FILE__ "NA.v"
`define __LINE__ 0
`define DVT_PATCH

// CONFIGURATION FILES (libmap) 
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/defines.sv"
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/class_1.sv"
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/class_2.sv"
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/class_3.sv"
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/class_4.sv"
`include "/home/student/akamien/dvt_predefined_projects_target/sv-GettingStarted/class_5.sv"
